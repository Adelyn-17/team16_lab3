module vga_char
