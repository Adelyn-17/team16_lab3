module vga_colorbar
