module vga_ctrl
