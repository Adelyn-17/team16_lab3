module vga_pic
