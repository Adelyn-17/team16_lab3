module vga_pic(
    input wire vga_clk,
    input wire sys_rst_n,
    input wire [9:0] pix_x,
    input wire [9:0] pix_y,

    output wire [15:0] pix_data  
);

parameter CHAR_B_H = 10'd192,  
          CHAR_B_V = 10'd208;  
			 
parameter CHAR_W = 10'd256,    
          CHAR_H = 10'd64;     
			 
parameter BLACK  = 16'h0000,   
          GOLDEN = 16'hFEC0;  

reg [255:0] char [63:0];  
wire [9:0] char_x;        
wire [9:0] char_y;        
reg [15:0] pix_data_reg;

assign char_x = ( (pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W))
                && (pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H)) )
                ? (pix_x - CHAR_B_H) : 10'd256; 

assign char_y = ( (pix_x >= CHAR_B_H) && (pix_x < (CHAR_B_H + CHAR_W))
                && (pix_y >= CHAR_B_V) && (pix_y < (CHAR_B_V + CHAR_H)) )
                ? (pix_y - CHAR_B_V) : 10'd64;   

assign pix_data = pix_data_reg;


initial begin
    char[0]  <= 256'h00000000000000000000000000000000;
    char[1]  <= 256'h00000000000000000000000000000000;
    char[2]  <= 256'h00000000000000000000000000000000;
    char[3]  <= 256'h00000000000000000000000000000000;
    char[4]  <= 256'h00000000000000000000000000000000;
    char[5]  <= 256'h00000000000000000000000000000000;
    char[6]  <= 256'h00000000000000000000000000000000;
    char[7]  <= 256'h00000000000000000000000000000000;
    char[8]  <= 256'h00000000000000000000000000000000;
    char[9]  <= 256'h00000000000000000000000000000000;
    char[10] <= 256'h00000000000000000000000000000000;
    char[11] <= 256'h00000000000000000000000000000000;
    char[12] <= 256'h00000000000000000000000000000000;
    char[13] <= 256'h00000000000000000000000000000000;
    char[14] <= 256'h00000000000000000000000000000000;
    char[15] <= 256'h00000000000000000000000000000000;
    char[16] <= 256'h00000000000000000000000000000000;
    char[17] <= 256'h00000000000000000000000000000000;
    char[18] <= 256'h00000000000000000000000000000000;
    char[19] <= 256'h00000000000000000000000000000000;
    char[20] <= 256'h00000000000000000000000000000000;
    char[21] <= 256'h00000000000000000000000000000000;
    char[22] <= 256'h00000000000000000000000000000000;
    char[23] <= 256'h00000000000000000000000000000000;
    char[24] <= 256'h00000000000000000000000000000000;
    char[25] <= 256'h00000000000000000000000000000000;
    char[26] <= 256'h000C3000000C30000003C000000FF000;
    char[27] <= 256'h000C3000000C30000007E000000FF000;
    char[28] <= 256'h000E7000000C3000000E700000018000;
    char[29] <= 256'h000E7000000C3000000E000000018000;
    char[30] <= 256'h000FF000000C30000007000000018000;
    char[31] <= 256'h000FF000000C30000003800000018000;
    char[32] <= 256'h000DB000000C30000000C00000018000;
    char[33] <= 256'h000DB000000C30000000600000018000;
    char[34] <= 256'h000C3000000C30000000700000018000;
    char[35] <= 256'h000C3000000E7000000E700000018000;
    char[36] <= 256'h000C30000007E0000007E00000018000;
    char[37] <= 256'h000C30000003C0000003C00000018000;
    char[38] <= 256'h00000000000000000000000000000000;
    char[39] <= 256'h00000000000000000000000000000000;
    char[40] <= 256'h00000000000000000000000000000000;
    char[41] <= 256'h00000000000000000000000000000000;
    char[42] <= 256'h00000000000000000000000000000000;
    char[43] <= 256'h00000000000000000000000000000000;
    char[44] <= 256'h00000000000000000000000000000000;
    char[45] <= 256'h00000000000000000000000000000000;
    char[46] <= 256'h00000000000000000000000000000000;
    char[47] <= 256'h00000000000000000000000000000000;
    char[48] <= 256'h00000000000000000000000000000000;
    char[49] <= 256'h00000000000000000000000000000000;
    char[50] <= 256'h00000000000000000000000000000000;
    char[51] <= 256'h00000000000000000000000000000000;
    char[52] <= 256'h00000000000000000000000000000000;
    char[53] <= 256'h00000000000000000000000000000000;
    char[54] <= 256'h00000000000000000000000000000000;
    char[55] <= 256'h00000000000000000000000000000000;
    char[56] <= 256'h00000000000000000000000000000000;
    char[57] <= 256'h00000000000000000000000000000000;
    char[58] <= 256'h00000000000000000000000000000000;
    char[59] <= 256'h00000000000000000000000000000000;
    char[60] <= 256'h00000000000000000000000000000000;
    char[61] <= 256'h00000000000000000000000000000000;
    char[62] <= 256'h00000000000000000000000000000000;
    char[63] <= 256'h00000000000000000000000000000000;
end


always @(posedge vga_clk or negedge sys_rst_n) begin
    if (sys_rst_n == 1'b0) begin
        pix_data_reg <= BLACK;
    end else if ( (char_x < CHAR_W) && (char_y < CHAR_H)  
                  && (char[char_y][char_x] == 1'b1) ) begin
        pix_data_reg <= GOLDEN;
    end else begin
        pix_data_reg <= BLACK;
    end
end

endmodule
